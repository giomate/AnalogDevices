// spin_sensor_receiver.v

// Generated using ACDS version 20.1 711

`timescale 1 ps / 1 ps
module spin_sensor_receiver (
		input  wire  clk_clk,       //   clk.clk
		input  wire  reset_reset_n  // reset.reset_n
	);

endmodule
