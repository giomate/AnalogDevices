-- spin_sensor_receiver_spin_sensor_receiver_0.vhd

-- Generated using ACDS version 20.1 711

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity spin_sensor_receiver_spin_sensor_receiver_0 is
	port (
		clk_clk       : in std_logic := '0'; --   clk.clk
		reset_reset_n : in std_logic := '0'  -- reset.reset_n
	);
end entity spin_sensor_receiver_spin_sensor_receiver_0;

architecture rtl of spin_sensor_receiver_spin_sensor_receiver_0 is
	component spin_sensor_receiver_spin_sensor_receiver_0_spin_sensor_receiver_0 is
	end component spin_sensor_receiver_spin_sensor_receiver_0_spin_sensor_receiver_0;

begin

	spin_sensor_receiver_0 : component spin_sensor_receiver_spin_sensor_receiver_0_spin_sensor_receiver_0
		port map (
		);

end architecture rtl; -- of spin_sensor_receiver_spin_sensor_receiver_0
